module add2(in,out);

input [7:0]in;
output [7:0]out;

assign out=in+2;

endmodule